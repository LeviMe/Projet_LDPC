
library ieee; 
use ieee.std_logic_1164.all;

-- Première tentative de réaliser l'encodeur LDPC du code CCSDS binaire 128, 256
-- encodage systématique: sortie = entrée & entrée x (partie droite de G)
-- produit scalaire avec chacune des lignes de la transposée, faite de la concaténation de 4 matrices circulantes.
-- Version 100% parralèle: l'ensemble du produit matriciel se fait en un seul cycle, sans process. 
-- Pas de signaux ajouté pour la synchronisation avec les autres modules. 
-- 1ere version pour évaluation première l'usage des ressources.
-- Préparé une version semi-série: pas de raison d'avoir un encodage aussi rapide si un appareil du meme type
-- fait le décodage avec nécessairement de multiples cycles d'horloges.

-- possible danger à utiliser les fonctions de décalage directement sur des vecteurs. https://stackoverflow.com/a/30556879
-- pas compilable ==> création de mes propres fonctions de décalage.

-- logique dupliquée avec des for dans des fonctions; Les for sont utilisables dans les fonctions ou les process seulement.
-- les deux limites du for sont incluses.

entity encoder is 

generic (
	constant K : integer := 128;
	constant N : integer := 256; 
	
	constant L0 :  std_logic_vector(127 downto 0):= x"7546f665fbf07eec75902581e7ebd072";
	constant L32 : std_logic_vector(127 downto 0):= x"c196638a4bfe987179a486f304419ca2";
	constant L64 : std_logic_vector(127 downto 0):= x"a1ecd4631cd81a9d8f0db2506ddad1d2";
	constant L96 : std_logic_vector(127 downto 0):= x"f5ea237904bd6e24b41212b8e73d62c5"
);

port (
	input :  in std_logic_vector(K-1 downto 0);
	output : out std_logic_vector(N-1 downto 0)
);

end encoder; 


architecture rtl of encoder is
 	function shift_circ_r(
		L: in std_logic_vector; index : in integer)
		return std_logic_vector is
		variable size: integer := L'Length;
		variable res : std_logic_vector(size-1 downto 0) := (others => '0');
		begin
			res := L(size-1-index downto 0) & L(size-1 downto size-index);
		return res;
		
	end function shift_circ_r;
	
	 function sum_xor (
		 in_vec    : in std_logic_vector)
		 return std_logic is
		 variable s : std_logic := '0';
		 begin
			 for i in in_vec'low to in_vec'high loop -- changé pour compiler valeur dans testbench. Attention: to -> croissant, dowto -> décroissant.
					s := s xor in_vec(i);
					--report std_logic'image(in_vec(i)) & std_logic'image(s) ;
			 end loop;
			 report "entree dans sum_xor" & std_logic'image(s);
		 return s;  
	  end function sum_xor;
	
	
	function circular_perm4(L : in std_logic_vector; index : in integer := 0)
	return  std_logic_vector is	
		variable  res : 	std_logic_vector(127 downto 0) := (others => '0');
		variable  mot :  	std_logic_vector(31  downto 0) := (others => '0');
		variable  mot_per :  	std_logic_vector(31  downto 0) := (others => '0');
		begin 
			decomp : for i in 0 to 3 loop
							mot := L((i+1)*32 -1 downto i*32); 
							mot_per := shift_circ_r(mot, index); 
							res((i+1)*32 - 1 downto i*32) := mot_per;
			end loop decomp;
			return res;
	end function;
	
	function encode(input: in std_logic_vector) return std_logic_vector is
		variable s_droite : std_logic_vector(127 downto 0) := (others => '0');
		begin
		for i in 0 to 31 loop
			s_droite(i) 	:=  sum_xor(input and circular_perm4(L0,  i));
			s_droite(i+32)  :=  sum_xor(input and circular_perm4(L32, i));
			s_droite(i+64)  :=  sum_xor(input and circular_perm4(L64, i));
			s_droite(i+96)  :=  sum_xor(input and circular_perm4(L96, i));
		end loop;
		
		return s_droite & input ;
	end function;

begin
	output <= encode(input);
end rtl;
